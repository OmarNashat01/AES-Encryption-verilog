module MixColumns(input data[127:0] byte, output reg[127:0] Sbyte);

always@()


endmodule

