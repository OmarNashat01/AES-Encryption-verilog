module AddRoundKey();

endmodule