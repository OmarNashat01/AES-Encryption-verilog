module MixColumns(input wire[127:0] byte, output reg[127:0] Sbyte);



endmodule

