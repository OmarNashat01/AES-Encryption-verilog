module LastRound(

						input wire[127:0] Keyin,
						input wire[127:0] Indata,
						
						output[127:0] data
						);
						
endmodule