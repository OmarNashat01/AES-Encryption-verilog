module KeyExpansion(
	input [3:0] round,
	input [31:0] keyin,
	output reg [31:0] keyout
);



endmodule